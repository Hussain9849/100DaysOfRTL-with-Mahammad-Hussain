module mux21(i0,i1,s,y);
   input i0,i1,s;
   output y;
   assign y = (s==1)?i1:i0;

endmodule
