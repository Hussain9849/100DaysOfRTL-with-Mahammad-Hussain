module Positive_d_latch(d,en,q,qb);
    input d,en;
	output q,qb;
	not n(w1,);
endmodule
