module SRlatch(S,R,Q,Qb);
   input S,R;
   output Q,Qb;
   wire Sb,Rb;
   nand g0(Q,Sb,Qb);
   nand g2(Qb,Rb,Q);
   nand g3(Sb,S,S);
   nand g4(Rb,R,R);
endmodule
