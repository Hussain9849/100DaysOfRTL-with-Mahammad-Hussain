module Mux_8_1(input [7:0] I,input [2:0] S,output Y);

  assign Y = (I[0] & ~S[2] & ~S[1] & ~S[0]) |
             (I[1] & ~S[2] & ~S[1] &  S[0]) |
             (I[2] & ~S[2] &  S[1] & ~S[0]) |
             (I[3] & ~S[2] &  S[1] &  S[0]) |
             (I[4] &  S[2] & ~S[1] & ~S[0]) |
             (I[5] &  S[2] & ~S[1] &  S[0]) |
             (I[6] &  S[2] &  S[1] & ~S[0]) |
             (I[7] &  S[2] &  S[1] &  S[0]);
endmodule

module Mux_8_1_TB;
  reg [7:0] I;
  reg [2:0] S;
  wire Y;

  Mux_8_1 UUT(.I(I), .S(S), .Y(Y));

  initial begin
    $display("Time\t  I       S2 S1 S0 | Y");
    $monitor("%g\t %b  %b  %b  %b | %b", $time,I, S[2], S[1], S[0], Y);

    // Test each input line
    I = 8'b00000001; S = 3'b000; #10;
    I = 8'b00000010; S = 3'b001; #10;
    I = 8'b00000100; S = 3'b010; #10;
    I = 8'b00001000; S = 3'b011; #10;
    I = 8'b00010000; S = 3'b100; #10;
    I = 8'b00100000; S = 3'b101; #10;
    I = 8'b01000000; S = 3'b110; #10;
    I = 8'b10000000; S = 3'b111; #10;
    $finish;
  end
endmodule

