module GrayToBinary_3bit(input g2, g1, g0, output b2, b1, b0);
  wire [3:0] I_b2;
  wire [3:0] I_b1;
  wire [3:0] I_b0;
  wire not_g0;
  not G2(not_g0, g0);
  assign I_b2 = {1'b1, 1'b1, 1'b0, 1'b0};                   
  assign I_b1 = {1'b0, 1'b1, 1'b1, 1'b0};                  
  assign I_b0 = {g0, not_g0, not_g0, g0};                   
  Mux_4_1 M1(.i(I_b2), .s1(g2), .s0(g1), .y(b2));
  Mux_4_1 M2(.i(I_b1), .s1(g2), .s0(g1), .y(b1));
  Mux_4_1 M3(.i(I_b0), .s1(g2), .s0(g1), .y(b0));
endmodule

module GrayToBinary_tb;
  reg g2, g1, g0;
  wire b2, b1, b0;
  GrayToBinary uut (.g2(g2), .g1(g1), .g0(g0),.b2(b2), .b1(b1), .b0(b0));
  initial begin
    $display("Time | g2 g1 g0 | b2 b1 b0");
    $monitor("%4t |  %b  %b  %b |  %b  %b  %b", $time, g2, g1, g0, b2, b1, b0);

    g2=0; g1=0; g0=0; #10;
    g2=0; g1=0; g0=1; #10;
    g2=0; g1=1; g0=0; #10;
    g2=0; g1=1; g0=1; #10;
    g2=1; g1=0; g0=0; #10;
    g2=1; g1=0; g0=1; #10;
    g2=1; g1=1; g0=0; #10;
    g2=1; g1=1; g0=1; #10;
    $finish;
  end
endmodule
