module Full_Sub_Using_8_1Mux(input A, B, Bin, output Diff, Borr);

  wire [2:0] Sel = {A, B, Bin};  // Sel = ABC
  wire [7:0] I_Diff = 8'b10010110;  
  wire [7:0] I_Borr = 8'b10001110;


  Mux_8_1 M1 (.Y(Diff), .S(Sel), .I(I_Diff));
  Mux_8_1 M2 (.Y(Borr), .S(Sel), .I(I_Borr));

endmodule

module Full_Sub_Using_8_1Mux_tb;

  reg A, B, Bin;
  wire Diff, Borr;

  Full_Sub_Using_8_1Mux uut (.A(A),.B(B),.Bin(Bin),.Diff(Diff),.Borr(Borr));

  initial begin
    $display("Time\t A B Bin |Diff Borr");
    $monitor("%g\t %b %b %b   | %b    %b", $time, A, B, Bin, Diff, Borr);

    A = 0; B = 0; Bin = 0; #10;
    A = 0; B = 0; Bin = 1; #10;
    A = 0; B = 1; Bin = 0; #10;
    A = 0; B = 1; Bin = 1; #10;
    A = 1; B = 0; Bin = 0; #10;
    A = 1; B = 0; Bin = 1; #10;
    A = 1; B = 1; Bin = 0; #10;
    A = 1; B = 1; Bin = 1; #10;

    $finish;
  end

endmodule

